// ************************************************ ******************** 
// >>>>>>>>>>>>>>>>>>>>>>>>> COPYRIGHT NOTICE < <<<<<<<<<<<<<<<<<<<<<<<< 
// ************************ ******************************************** 
// File name: divide_tb .v 
// Module name: divide_tb 
// Author: STEP 
// Description: clock divider 
// Web: www.stepfpga.com 
// 
// ------------------ -------------------------------------------------- 
// Code Revision History: 
// ------------------------------------------ -------------------------- 
// Version: |Mod. Date: |Changes Made:
// V1.0 |2017/03/02 |Initial ver
// ------------------------------------------------ -------------------- 
// Module Function: divide.v test file of clock divider

`timescale 1ns / 100ps   //simulation time unit/time accuracy, the time unit must be greater than or equal to the time accuracy

module divide_tb ();  //The test file is also a module, because it is used for simulation, there is no need for input and output signals
	
	reg clk, rst_n;   //The definition of the excitation signal that needs to be generated, the excitation signal needs to be generated by the process block, so it is defined as a reg type variable 
	wire clkout;      //The output signal definition that needs to be observed is defined as a wire type variable
	
	// Initialization process block
	initial
	begin
		clk = 0;
		rst_n = 0;
		# 25
		rst_n = 1;	
	end
	
	always #10 clk = ~clk;  //Invert the clk signal every 10ns, that is, generate a clk with a clock cycle of 20ns, and the frequency is 50MHz  
		
		divide #(.WIDTH(4), .N(11)) u1(   //#The following () is for parameter passing, if no parameter is passed, it is the default value of the parameter in the called module 
                                            // divide represents a desired embodiment of the module name, the name U1 is the embodiment of our definition, must begin with a letter 
		            .clk(clk),             // O signal name represents a signal connection module itself .clk defined;. (clk) represents here we define the excitation signal
					.rst_n(rst_n),         // different ports signal name // defined in the testbench and can be invoked in the module
				    .clkout(CLKOUT)
					);

endmodule